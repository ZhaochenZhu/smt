VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
CLEARANCEMEASURE EUCLIDEAN ;

MACRO INVx1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx1_ASAP7_75t_R 0 0 ;
  SIZE 0.084 BY 0.216 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.105 0.072 0.147 0.192 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.273 0.072 0.315 0.192 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.000 0.192 0.084 0.240 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.000 -0.024 0.084 0.024 ;
    END
  END VSS
END INVx1_ASAP7_75t_R

SITE coreSite
	CLASS CORE ;
	SYMMETRY X Y R90 ;
	SIZE 0.084 BY 0.216 ;
END coreSite

END LIBRARY
