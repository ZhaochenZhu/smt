VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
CLEARANCEMEASURE EUCLIDEAN ;

SITE coreSite
	CLASS CORE ;
	SYMMETRY X Y R90 ;
	SIZE 0.084 BY 0.0 ;
END coreSite

END LIBRARY
